LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY ALU IS
	GENERIC (m:integer:=16);
	PORT(a,b: IN STD_LOGIC_VECTOR(m-1 DOWNTO 0);
        s : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        flagsIn : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        c : OUT STD_LOGIC_VECTOR(m-1 DOWNTO 0)
        flagsOut: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)); -- C - N - Z
END ENTITY ALU;

ARCHITECTURE ALUArch OF ALU IS

BEGIN


END ARCHITECTURE;

