LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY MUX2x1 IS
	GENERIC (n:INTEGER:=16);
	PORT(a,b: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		s : IN STD_LOGIC;
		c : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0));
END ENTITY MUX2x1;

ARCHITECTURE MUX2x1Arch OF MUX2x1 IS

BEGIN

c <= a WHEN s = '0' 
ELSE b WHEN s = '1';

END ARCHITECTURE;
