LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY DataHazard IS
    port()
END ENTITY DataHazard;

Architecture DataHazardArch OF DataHazard

begin


END Architecture