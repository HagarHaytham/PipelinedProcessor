ENTITY fetchControl IS
	PORT(	
